----------------------------------------------------------------------------
----------------------------------------------------------------------------
--
-- Copyright 2016,2017 International Business Machines
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions AND
-- limitations under the License.
--
----------------------------------------------------------------------------
----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity action_axi_slave is
	generic (
		-- Users to add parameters here

		-- User parameters ends
		-- Do not modify the parameters beyond this line

		-- Width of S_AXI data bus
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		-- Width of S_AXI address bus
		C_S_AXI_ADDR_WIDTH	: integer	:= 6
	);
	port (
		-- Users to add ports here
                reg_0x10_i      : in  std_logic_vector(31 downto 0);
                reg_0x14_i      : in  std_logic_vector(31 downto 0);
                reg_0x20_o      : out std_logic_vector(31 downto 0);
                reg_0x30_o      : out std_logic_vector(31 downto 0);
                reg_0x34_o      : out std_logic_vector(31 downto 0);
                reg_0x38_o      : out std_logic_vector(31 downto 0);
                reg_0x3c_o      : out std_logic_vector(31 downto 0);
                reg_0x40_o      : out std_logic_vector(31 downto 0);
                reg_0x44_o      : out std_logic_vector(31 downto 0);
				reg_0x48_o      : out std_logic_vector(31 downto 0);
                int_enable_o    : out std_logic;
                app_start_o     : out std_logic;
                app_done_i      : in  std_logic;
                app_ready_i     : in  std_logic;
                app_idle_i      : in  std_logic;

        -- for debug only
                after_done_i                : in std_logic;
                after_all_wr_ack_i          : in std_logic;
                after_rd_done_i             : in std_logic;
                after_first_wr_ack_i        : in std_logic;
                after_wr_data_sent_i        : in std_logic;
                after_first_wr_rqt_ack_i    : in std_logic;
                after_first_wr_rqt_i        : in std_logic;
                after_start_i               : in std_logic;
                after_first_wr_ready_i      : in std_logic;
                after_first_wr_valid_i      : in std_logic;
                process_cnt_i               : in std_logic_vector(25 downto 0);
                

        -- Registers from 0x60 to 0x7c are reserved for the debug in this application 

                --reg_0x60_i      : in std_logic_vector(31 downto 0);
                --reg_0x64_i      : in std_logic_vector(31 downto 0);
                --reg_0x68_i      : in std_logic_vector(31 downto 0);
                --reg_0x6c_i      : in std_logic_vector(31 downto 0);
                --reg_0x70_i      : in std_logic_vector(31 downto 0);
                --reg_0x74_i      : in std_logic_vector(31 downto 0);
                --reg_0x78_i      : in std_logic_vector(31 downto 0);
                --reg_0x7c_i      : in std_logic_vector(31 downto 0);
               
                
		-- User ports ends
		-- Do not modify the ports beyond this line

		-- Global Clock Signal
		S_AXI_ACLK	: in std_logic;
		-- Global Reset Signal. This Signal is Active LOW
		S_AXI_ARESETN	: in std_logic;
		-- Write address (issued by master, acceped by Slave)
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
--		-- Write channel Protection type. This signal indicates the
--    		-- privilege and security level of the transaction, and whether
--    		-- the transaction is a data access or an instruction access.
--		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		-- Write address valid. This signal indicates that the master signaling
    		-- valid write address and control information.
		S_AXI_AWVALID	: in std_logic;
		-- Write address ready. This signal indicates that the slave is ready
    		-- to accept an address and associated control signals.
		S_AXI_AWREADY	: out std_logic;
		-- Write data (issued by master, acceped by Slave) 
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Write strobes. This signal indicates which byte lanes hold
    		-- valid data. There is one write strobe bit for each eight
    		-- bits of the write data bus.    
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		-- Write valid. This signal indicates that valid write
    		-- data and strobes are available.
		S_AXI_WVALID	: in std_logic;
		-- Write ready. This signal indicates that the slave
    		-- can accept the write data.
		S_AXI_WREADY	: out std_logic;
		-- Write response. This signal indicates the status
    		-- of the write transaction.
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		-- Write response valid. This signal indicates that the channel
    		-- is signaling a valid write response.
		S_AXI_BVALID	: out std_logic;
		-- Response ready. This signal indicates that the master
    		-- can accept a write response.
		S_AXI_BREADY	: in std_logic;
		-- Read address (issued by master, acceped by Slave)
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
--		-- Protection type. This signal indicates the privilege
--    		-- and security level of the transaction, and whether the
--    		-- transaction is a data access or an instruction access.
--		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		-- Read address valid. This signal indicates that the channel
    		-- is signaling valid read address and control information.
		S_AXI_ARVALID	: in std_logic;
		-- Read address ready. This signal indicates that the slave is
    		-- ready to accept an address and associated control signals.
		S_AXI_ARREADY	: out std_logic;
		-- Read data (issued by slave)
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		-- Read response. This signal indicates the status of the
    		-- read transfer.
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		-- Read valid. This signal indicates that the channel is
    		-- signaling the required read data.
		S_AXI_RVALID	: out std_logic;
		-- Read ready. This signal indicates that the master can
    		-- accept the read data and response information.
		S_AXI_RREADY	: in std_logic
	);
end action_axi_slave;

architecture action_axi_slave of action_axi_slave is

	-- AXI4LITE signals
	signal axi_awaddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_awready	: std_logic;
	signal axi_wready	: std_logic;
	signal axi_bresp	: std_logic_vector(1 downto 0);
	signal axi_bvalid	: std_logic;
	signal axi_araddr	: std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
	signal axi_arready	: std_logic;
	signal axi_rdata	: std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal axi_rresp	: std_logic_vector(1 downto 0);
	signal axi_rvalid	: std_logic;

	-- Example-specific design signals
	-- local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	-- ADDR_LSB is used for addressing 32/64 bit registers/memories
	-- ADDR_LSB = 2 for 32 bits (n downto 2)
	-- ADDR_LSB = 3 for 64 bits (n downto 3)
	constant ADDR_LSB          : integer := (C_S_AXI_DATA_WIDTH/32)+ 1;
	constant OPT_MEM_ADDR_BITS : integer := 5;
	------------------------------------------------
	---- Signals for user logic register space example
	--------------------------------------------------
	---- Number of Slave Registers 16
	signal slv_reg0	        : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg0_new     : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg1         : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg2         : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg3         : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg8         : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg12	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg13	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg14	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg15	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg16	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg17	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg18	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg19	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg_rden	    : std_logic;
	signal slv_reg_wren	    : std_logic;
	signal reg_data_out	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal byte_index	    : integer;
    
    signal idle_q           : std_logic;
    signal app_start_q      : std_logic;
    signal app_done_q       : std_logic;
    signal slv_reg0_bit0_q  : std_logic;

-- for debugging only
	signal slv_reg24	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg25	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg26	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg27	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg28	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg29	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg30	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal slv_reg31	    : std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
	signal after_done_q             : std_logic;
	signal after_all_wr_ack_q       : std_logic;
	signal after_rd_done_q          : std_logic;
	signal after_first_wr_ack_q     : std_logic;
	signal after_wr_data_sent_q     : std_logic;
	signal after_first_wr_rqt_ack_q : std_logic;
	signal after_first_wr_rqt_q     : std_logic;
	signal after_start_q            : std_logic;
    signal after_first_wr_ready_q   : std_logic;
    signal after_first_wr_valid_q   : std_logic;
    signal process_cnt_q            : std_logic_vector(25 downto 0);

begin
	-- I/O Connections assignments

    int_enable_o    <= slv_reg1(0);
	S_AXI_AWREADY	<= axi_awready;
	S_AXI_WREADY	<= axi_wready;
	S_AXI_BRESP	<= axi_bresp;
	S_AXI_BVALID	<= axi_bvalid;
	S_AXI_ARREADY	<= axi_arready;
	S_AXI_RDATA	<= axi_rdata;
	S_AXI_RRESP	<= axi_rresp;
	S_AXI_RVALID	<= axi_rvalid;
	-- Implement axi_awready generation
	-- axi_awready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
	-- de-asserted when reset is low.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awready <= '0';
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1') then
	        -- slave is ready to accept write address when
	        -- there is a valid write address and write data
	        -- on the write address and data bus. This design 
	        -- expects no outstanding transactions. 
	        axi_awready <= '1';
	      else
	        axi_awready <= '0';
	      end if;
	    end if;
	  end if;
	end process;

	-- Implement axi_awaddr latching
	-- This process is used to latch the address when both 
	-- S_AXI_AWVALID and S_AXI_WVALID are valid. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_awaddr <= (others => '0');
	    else
	      if (axi_awready = '0' and S_AXI_AWVALID = '1' and S_AXI_WVALID = '1') then
	        -- Write Address latching
	        axi_awaddr <= S_AXI_AWADDR;
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_wready generation
	-- axi_wready is asserted for one S_AXI_ACLK clock cycle when both
	-- S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
	-- de-asserted when reset is low. 

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_wready <= '0';
	    else
	      if (axi_wready = '0' and S_AXI_WVALID = '1' and S_AXI_AWVALID = '1') then
	          -- slave is ready to accept write data when 
	          -- there is a valid write address and write data
	          -- on the write address and data bus. This design 
	          -- expects no outstanding transactions.           
	          axi_wready <= '1';
	      else
	        axi_wready <= '0';
	      end if;
	    end if;
	  end if;
	end process; 

	-- Implement memory mapped register select and write logic generation
	-- The write data is accepted and written to memory mapped registers when
	-- axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
	-- select byte enables of slave registers while writing.
	-- These registers are cleared when reset (active low) is applied.
	-- Slave register write enable is asserted when valid address and data are available
	-- and the slave is ready to accept the write address and write data.
	slv_reg_wren <= axi_wready and S_AXI_WVALID and axi_awready and S_AXI_AWVALID ;

	process (S_AXI_ACLK)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS-1 downto 0); 
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      slv_reg0 <= (others => '0');
	      slv_reg1 <= (others => '0');
	      slv_reg2 <= (others => '0');
	      slv_reg3 <= (others => '0');
	      slv_reg8 <= (others => '0');
	      slv_reg12 <= (others => '0');
	      slv_reg13 <= (others => '0');
	      slv_reg14 <= (others => '0');
	      slv_reg15 <= (others => '0');
	      slv_reg16 <= (others => '0');
	      slv_reg17 <= (others => '0');
	      slv_reg18 <= (others => '0');
	      slv_reg19 <= (others => '0');
	    else
	      loc_addr := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS-1 downto ADDR_LSB);
	      if (slv_reg_wren = '1') then
	        case loc_addr is
	          when b"00000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 0
	                slv_reg0(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00001" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 1
	                slv_reg1(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00010" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 2
	                slv_reg2(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"00011" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 3
	                slv_reg3(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 8
	                slv_reg8(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01100" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 12
	                slv_reg12(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01101" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 13
	                slv_reg13(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01110" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 14
	                slv_reg14(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"01111" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 15
	                slv_reg15(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10000" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 16
	                slv_reg16(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10001" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 17
	                slv_reg17(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10010" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 18
	                slv_reg18(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;
	          when b"10011" =>
	            for byte_index in 0 to (C_S_AXI_DATA_WIDTH/8-1) loop
	              if ( S_AXI_WSTRB(byte_index) = '1' ) then
	                -- Respective byte enables are asserted as per write strobes                   
	                -- slave registor 19
	                slv_reg19(byte_index*8+7 downto byte_index*8) <= S_AXI_WDATA(byte_index*8+7 downto byte_index*8);
	              end if;
	            end loop;

	          when others =>
	            slv_reg0 <= slv_reg0;
	            slv_reg1 <= slv_reg1;
	            slv_reg2 <= slv_reg2;
	            slv_reg3 <= slv_reg3;
	            slv_reg8 <= slv_reg8;
	            slv_reg12 <= slv_reg12;
	            slv_reg13 <= slv_reg13;
	            slv_reg14 <= slv_reg14;
	            slv_reg15 <= slv_reg15;
	            slv_reg16 <= slv_reg16;
	            slv_reg17 <= slv_reg17;
	            slv_reg18 <= slv_reg18;
	            slv_reg19 <= slv_reg19;
	        end case;
	      end if;
              if app_start_q = '1' then
                slv_reg0(0) <= '0';
              end if;  
	    end if;
	  end if;                   
	end process; 

	-- Implement write response logic generation
	-- The write response and response valid signals are asserted by the slave 
	-- when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
	-- This marks the acceptance of address and indicates the status of 
	-- write transaction.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_bvalid  <= '0';
	      axi_bresp   <= "00"; --need to work more on the responses
	    else
	      if (axi_awready = '1' and S_AXI_AWVALID = '1' and axi_wready = '1' and S_AXI_WVALID = '1' and axi_bvalid = '0'  ) then
	        axi_bvalid <= '1';
	        axi_bresp  <= "00"; 
	      elsif (S_AXI_BREADY = '1' and axi_bvalid = '1') then   --check if bready is asserted while bvalid is high)
	        axi_bvalid <= '0';                                 -- (there is a possibility that bready is always asserted high)
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arready generation
	-- axi_arready is asserted for one S_AXI_ACLK clock cycle when
	-- S_AXI_ARVALID is asserted. axi_awready is 
	-- de-asserted when reset (active low) is asserted. 
	-- The read address is also latched when S_AXI_ARVALID is 
	-- asserted. axi_araddr is reset to zero on reset assertion.

	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then 
	    if S_AXI_ARESETN = '0' then
	      axi_arready <= '0';
	      axi_araddr  <= (others => '1');
	    else
	      if (axi_arready = '0' and S_AXI_ARVALID = '1') then
	        -- indicates that the slave has acceped the valid read address
	        axi_arready <= '1';
	        -- Read Address latching 
	        axi_araddr  <= S_AXI_ARADDR;           
	      else
	        axi_arready <= '0';
	      end if;
	    end if;
	  end if;                   
	end process; 

	-- Implement axi_arvalid generation
	-- axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
	-- S_AXI_ARVALID and axi_arready are asserted. The slave registers 
	-- data are available on the axi_rdata bus at this instance. The 
	-- assertion of axi_rvalid marks the validity of read data on the 
	-- bus and axi_rresp indicates the status of read transaction.axi_rvalid 
	-- is deasserted on reset (active low). axi_rresp and axi_rdata are 
	-- cleared to zero on reset (active low).  
	process (S_AXI_ACLK)
	begin
	  if rising_edge(S_AXI_ACLK) then
	    if S_AXI_ARESETN = '0' then
	      axi_rvalid <= '0';
	      axi_rresp  <= "00";
	    else
	      if (axi_arready = '1' and S_AXI_ARVALID = '1' and axi_rvalid = '0') then
	        -- Valid read data is available at the read data bus
	        axi_rvalid <= '1';
	        axi_rresp  <= "00"; -- 'OKAY' response
	      elsif (axi_rvalid = '1' and S_AXI_RREADY = '1') then
	        -- Read data is accepted by the master
	        axi_rvalid <= '0';
	      end if;            
	    end if;
	  end if;
	end process;

	-- Implement memory mapped register select and read logic generation
	-- Slave register read enable is asserted when valid address is available
	-- and the slave is ready to accept the read address.
	slv_reg_rden <= axi_arready and S_AXI_ARVALID and (not axi_rvalid) ;

	process (slv_reg0_new, slv_reg1, slv_reg2, slv_reg3, reg_0x10_i, reg_0x14_i, slv_reg8, slv_reg12, slv_reg13, slv_reg14, slv_reg15, slv_reg16, slv_reg17, slv_reg18, slv_reg19, axi_araddr)
	variable loc_addr :std_logic_vector(OPT_MEM_ADDR_BITS-1 downto 0);
	begin
	    -- Address decoding for reading registers
	    loc_addr := axi_araddr(ADDR_LSB + OPT_MEM_ADDR_BITS-1 downto ADDR_LSB);
	    case loc_addr is
	      when b"00000" =>
	        reg_data_out <= slv_reg0_new;  -- 0x00
	      when b"00001" =>
	        reg_data_out <= slv_reg1;      -- 0x04
	      when b"00010" =>
	        reg_data_out <= slv_reg2;      -- 0x08
	      when b"00011" =>
	        reg_data_out <= slv_reg3;      -- 0x0c
	      when b"00100" =>
	        reg_data_out <= reg_0x10_i;    -- 0x10    
	      when b"00101" =>
	        reg_data_out <= reg_0x14_i;    -- 0x14
	      when b"01000" =>                  
	        reg_data_out <= slv_reg8;      -- 0x20
	      when b"01100" =>                  
	        reg_data_out <= slv_reg12;     -- 0x30
	      when b"01101" =>                  
	        reg_data_out <= slv_reg13;     -- 0x34
	      when b"01110" =>                  
	        reg_data_out <= slv_reg14;     -- 0x38
	      when b"01111" =>                  
	        reg_data_out <= slv_reg15;     -- 0x3c
	      when b"10000" =>                  
	        reg_data_out <= slv_reg16;     -- 0x40
	      when b"10001" =>                  
	        reg_data_out <= slv_reg17;     -- 0x44
	      when b"10010" =>                  
	        reg_data_out <= slv_reg18;     -- 0x48
	      when b"10011" =>                  
	        reg_data_out <= slv_reg19;     -- 0x4c
          -- the following registers are read-only for debugging in this application
          when b"11000" =>
            reg_data_out <= slv_reg24;     -- 0x60
          when b"11001" =>
            reg_data_out <= slv_reg25;     -- 0x64
          when b"11010" =>
            reg_data_out <= slv_reg26;     -- 0x68
          when b"11011" =>
            reg_data_out <= slv_reg27;     -- 0x6c
          when b"11100" =>
            reg_data_out <= slv_reg28;     -- 0x70
          when b"11101" =>
            reg_data_out <= slv_reg29;     -- 0x74
          when b"11110" =>
            reg_data_out <= slv_reg30;     -- 0x78
          when b"11111" =>
            reg_data_out <= slv_reg31;     -- 0x7c

	      when others =>
	        reg_data_out  <= (others => '0');
	    end case;
	end process;

    -- Debugging Register
--    slv_reg24 <= (others=>'0');
--    slv_reg25 <= (others=>'0');
    slv_reg26 <= (others=>'0');
    slv_reg27 <= (others=>'0');
    slv_reg28 <= (others=>'0');
    slv_reg29 <= (others=>'0');
    slv_reg30 <= (others=>'0');
    slv_reg31 <= (others=>'0');

    slv_reg25   <= slv_reg31(31 downto 26) & process_cnt_q(25 downto 0);

    -- after_df_valid_q & after_first_data_read_q 
    -- after_first_rd_ready_q & after_first_rd_valid_q & after_done_q & after_all_wr_ack_q 
    -- after_rd_done_q & after_first_wr_ack_q & after_wr_data_sent_q & after_first_wr_ready_q
    -- after_first_wr_valid_q & after_first_wr_rqt_ack_q & after_first_wr_rqt_q & after_start_q 
    -- app_ready_i & idle_q & app_done_q & app_start_q;
    slv_reg24 <= slv_reg28(31 downto 14) & after_done_q & after_all_wr_ack_q & after_rd_done_q & after_first_wr_ack_q & after_wr_data_sent_q & after_first_wr_ready_q & after_first_wr_valid_q & after_first_wr_rqt_ack_q & after_first_wr_rqt_q & after_start_q & app_ready_i & idle_q & app_done_q & app_start_q;
    

	process( S_AXI_ACLK ) is
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
            after_done_q                <= '0';
            after_all_wr_ack_q          <= '0';
            after_rd_done_q             <= '0';
            after_first_wr_ack_q        <= '0';
            after_wr_data_sent_q        <= '0';
            after_first_wr_rqt_ack_q    <= '0';
            after_first_wr_rqt_q        <= '0';
            after_start_q               <= '0';
            after_first_wr_ready_q      <= '0';
            after_first_wr_valid_q      <= '0';
            process_cnt_q               <= (others=>'0');
	    else
            after_done_q                <= after_done_i;
            after_all_wr_ack_q          <= after_all_wr_ack_i;
            after_rd_done_q             <= after_rd_done_i;
            after_first_wr_ack_q        <= after_first_wr_ack_i;
            after_wr_data_sent_q        <= after_wr_data_sent_i;
            after_first_wr_rqt_ack_q    <= after_first_wr_rqt_ack_i;
            after_first_wr_rqt_q        <= after_first_wr_rqt_i;
            after_start_q               <= after_start_i;
            after_first_wr_ready_q      <= after_first_wr_ready_i;
            after_first_wr_valid_q      <= after_first_wr_valid_i;
            process_cnt_q               <= process_cnt_i;
	    end if;
	  end if;
	end process;

	-- Output register or memory read data
	process( S_AXI_ACLK ) is
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	      axi_rdata  <= (others => '0');
	    else
	      if (slv_reg_rden = '1') then
	        -- When there is a valid read address (S_AXI_ARVALID) with 
	        -- acceptance of read address by the slave (axi_arready), 
	        -- output the read dada 
	        -- Read address mux
	          axi_rdata <= reg_data_out;     -- register read data
	      end if;   
	    end if;
	  end if;
	end process;

        
        
	-- Add user logic here
        -- Reiner

        app_start_o     <= app_start_q;
        reg_0x20_o      <= slv_reg8;
        reg_0x30_o      <= slv_reg12;
        reg_0x34_o      <= slv_reg13;
        reg_0x38_o      <= slv_reg14;
        reg_0x3c_o      <= slv_reg15;
        reg_0x40_o      <= slv_reg16;
        reg_0x44_o      <= slv_reg17;
		reg_0x48_o		<= slv_reg18;
        process( S_AXI_ACLK ) is
          variable app_done_i_q    : std_logic;
          
          variable loc_addr        :std_logic_vector(OPT_MEM_ADDR_BITS-1 downto 0); 
	begin
	  if (rising_edge (S_AXI_ACLK)) then
	    if ( S_AXI_ARESETN = '0' ) then
	      app_start_q     <=    '0';
	      app_done_q      <=    '0';
              app_done_i_q    :=    '0';
              slv_reg0_bit0_q <=    '0';
              idle_q          <=    '0';
     	    else
              idle_q          <= app_idle_i;
              slv_reg0_bit0_q <= slv_reg0(0);
              app_done_i_q    := app_done_i;
              loc_addr        := axi_awaddr(ADDR_LSB + OPT_MEM_ADDR_BITS-1 downto ADDR_LSB);
              -- clear ap_done bit when register is read
              if slv_reg_rden = '1'and loc_addr = "00000"  then
                app_done_q     <= '0';
              end if;  
	      if (app_done_i_q = '0' and app_done_i = '1') then
                app_done_q     <= '1';
	      end if;
              if slv_reg0_bit0_q = '0' and slv_reg0(0) = '1' then
                app_start_q <= '1';
              end if;
              if idle_q = '1' and app_idle_i = '0' then
                app_start_q <= '0';
              end if;
                
	    end if;
	  end if;
	end process;
        slv_reg0_new <= slv_reg0 (31 downto 4) & app_ready_i & idle_q & app_done_q & app_start_q ;

        
	-- User logic ends

end action_axi_slave;
